library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mux is
--  Port ( );
end mux;

architecture Behavioral of mux is

begin


end Behavioral;
