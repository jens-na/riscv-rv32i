library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity pc is
--  Port ( );
end pc;

architecture Behavioral of pc is



begin


end Behavioral;
