library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

use work.utils.all;
use work.opcodes.all;
use work.interfaces.all;

entity main is
  Port (
    clk: in std_logic
  );
end main;

architecture Behavioral of main is
begin

end Behavioral;