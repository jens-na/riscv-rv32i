library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity registerfile is
--  Port ( );
end registerfile;

architecture Behavioral of registerfile is

begin


end Behavioral;
